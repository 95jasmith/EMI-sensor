module Toggle_Pin_Test
	(output i_Tx_On,
	 input SS);
	 
	 assign i_Tx_On = SS;
	 
endmodule